`ifndef ALIGNER_ENV_PKG
	`define ALIGNER_ENV_PKG

//`include "uvm_macros.svh" 

package aligner_env_pkg; 
	import uvm_pkg::*; 

`include "aligner_env.sv" 

endpackage

`endif