`ifndef APB_TYPES
	`define APB_TYPES


typedef virtual apb_interface apb_virtual_interface; 


`endif